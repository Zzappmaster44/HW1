`timescale 1ns/1ns
module adder(sum, cOut, A, B, cIn);
  
  output  sum, cOut;
  input   A, B, cIn;
  
  wire w1,w2,w3;
  
  xor #20 g1 (w1,A,B);
  xor #20 g2 (sum,w1,cIn);
  
  and #10 g3 (w2,w1,cIn);
  and #10 g4 (w3,A,B);
  
  or  #10 g5 (cOut,w2,w3);
  
endmodule
