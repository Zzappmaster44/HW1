library verilog;
use verilog.vl_types.all;
entity testBench_B is
end testBench_B;
