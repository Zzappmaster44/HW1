library verilog;
use verilog.vl_types.all;
entity testBench_S is
end testBench_S;
