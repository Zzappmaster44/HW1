library verilog;
use verilog.vl_types.all;
entity prob6_structual is
    port(
        \OUT\           : out    vl_logic;
        E               : in     vl_logic;
        W               : in     vl_logic;
        clk             : in     vl_logic
    );
end prob6_structual;
