library verilog;
use verilog.vl_types.all;
entity testBench is
end testBench;
